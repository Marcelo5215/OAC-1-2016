library	ieee;
use	ieee.std_logic_1164.all;
use	ieee.numeric_std.all;
use	ieee.math_real.all;
USE IEEE.numeric_std.ALL;

entity testbench_REG_BANK is
	generic(  DATA_WIDTH    : natural := 32;
		  ADDRESS_WIDTH : natural := 5 );
end testbench_REG_BANK;

architecture testbench_REG_BANK_arch of testbench_REG_BANK is

    component REG_BANK

    	generic(  DATA_WIDTH    : natural := 32;
		  ADDRESS_WIDTH : natural := 5 );

    	port (  clk, wren           : in std_logic;
		radd1, radd2, wadd  : in std_logic_vector(ADDRESS_WIDTH - 1 downto 0);
		wdata               : in std_logic_vector(DATA_WIDTH    - 1 downto 0);
		rdata1, rdata2      : out std_logic_vector(DATA_WIDTH   - 1 downto 0));

    end component;

     --Inputs
    signal clk   : std_logic;
    signal wren  : std_logic;
    signal radd1 : std_logic_vector(ADDRESS_WIDTH-1 downto 0) := (others => '0');
    signal radd2 : std_logic_vector(ADDRESS_WIDTH-1 downto 0) := (others => '0');
    signal wadd  : std_logic_vector(ADDRESS_WIDTH-1 downto 0) := (others => '0');
    signal wdata : std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');

    --Outputs
    signal rdata1 : std_logic_vector(DATA_WIDTH-1 downto 0);
    signal rdata2 : std_logic_vector(DATA_WIDTH-1 downto 0);

begin


    utt: REG_BANK port map (
        clk => clk,
        wren => wren,
        radd1 => radd1,
        radd2 => radd2,
        wadd => wadd,
        wdata => wdata,
        rdata1 => rdata1,
        rdata2 => rdata2
    );



    test : process
    begin

		--Teste escrita e leitura reg(1)
		wadd <= (0 => '1', 1 => '0', 2 => '0', 3 => '0', 4 => '0');
		wdata <= (0 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		--Apenas radd1
		radd1 <= (0 => '1',others => '0');
		radd2 <= (others => '0');
		wait for 100 ns;
		
		--Apenas radd2
		radd1 <= (others => '0');
		radd2 <= (0 => '1',others => '0');
		wait for 100 ns;

		--Ambos radd
		radd1 <= (0 => '1',others => '0');
		radd2 <= (0 => '1',others => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(2)
		wadd <= (0 => '0', 1 => '1', 2 => '0', 3 => '0', 4 => '0');
		wdata <= (0 => '1', 1 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', others => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '1', others => '0');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', others => '0');
		radd2 <= (0 => '0', 1 => '1', others => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(3)
		wadd <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', others => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '1', others => '0');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', others => '0');
		radd2 <= (0 => '1', 1 => '1', others => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(4)
		wadd <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(5)
		wadd <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '0');
		wait for 100 ns;


		--Teste escrita e leitura reg(6)
		wadd <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		wait for 100 ns;


		--Teste escrita e leitura reg(7)
		wadd <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '0');
		wait for 100 ns;


		--Teste escrita e leitura reg(8)
		wadd <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(9)
		wadd <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1', 8 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (00 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(10)
		wadd <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1', 8 => '1', 9 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(11)
		wadd <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1', 8 => '1',
		9 => '1', 10 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(12)
		wadd <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(13)
		wadd <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(14)
		wadd <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(15)
		wadd <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '0');
		wait for 100 ns;

		--Teste escrita e leitura reg(16)
		wadd <= (0 => '0', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		radd2 <= (0 => '0', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(17)
		wadd <= (0 => '1', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		radd2 <= (0 => '1', 1 => '0', 2 => '0', 3 => '0', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(18)
		wadd <= (0 => '0', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		radd2 <= (0 => '0', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(19)
		wadd <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		radd2 <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(20)
		wadd <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		radd2 <= (0 => '0', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(21)
		wadd <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		radd2 <= (0 => '1', 1 => '0', 2 => '1', 3 => '0', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(22)
		wadd <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		radd2 <= (0 => '0', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(23)
		wadd <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		radd2 <= (0 => '1', 1 => '1', 2 => '1', 3 => '0', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(24)
		wadd <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', 23 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		radd2 <= (0 => '0', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(25)
		wadd <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', 23 => '1',
		24 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		radd2 <= (0 => '1', 1 => '0', 2 => '0', 3 => '1', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(26)
		wadd <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', 23 => '1',
		24 => '1', 25 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		radd2 <= (0 => '0', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(27)
		wadd <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', 23 => '1',
		24 => '1', 25 => '1', 26 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		radd2 <= (0 => '1', 1 => '1', 2 => '0', 3 => '1', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(28)
		wadd <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', 23 => '1',
		24 => '1', 25 => '1', 26 => '1', 27 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		radd2 <= (0 => '0', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(29)
		wadd <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', 23 => '1',
		24 => '1', 25 => '1', 26 => '1', 27 => '1', 28 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		radd2 <= (0 => '1', 1 => '0', 2 => '1', 3 => '1', 4 => '1');
		wait for 100 ns;


		--Teste escrita e leitura reg(30)
		wadd <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', 23 => '1',
		24 => '1', 25 => '1', 26 => '1', 27 => '1', 28 => '1', 29 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		radd2 <= (0 => '0', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		wait for 100 ns;

		--Teste escrita e leitura reg(31)
		wadd <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		wdata <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1', 5 => '1', 6 => '1', 7 => '1',
		8 => '1', 9 => '1', 10 => '1', 11 => '1', 12 => '1', 13 => '1', 14 => '1', 15 => '1',
		16 => '1', 17 => '1', 18 => '1', 19 => '1', 20 => '1', 21 => '1', 22 => '1', 23 => '1',
		24 => '1', 25 => '1', 26 => '1', 27 => '1', 28 => '1', 29 => '1', 30 => '1', others => '0');
		wren <= '1';
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		radd2 <= (others => '0');
		wait for 100 ns;

		radd1 <= (others => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		wait for 100 ns;

		radd1 <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		radd2 <= (0 => '1', 1 => '1', 2 => '1', 3 => '1', 4 => '1');
		wait for 100 ns;

		-- Teste reg(0)
		wadd <= (0 => '0', 1 => '0', 2 => '0', 3 => '0', 4 => '0');
		wdata <= (others => '1');
		wren <= '1';
		radd1 <= (others => '0');
		wait for 100 ns;

		--Leitura e escrita no mesmo ciclo
		wadd <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '0');
		wdata <= (others => '1');
		wren <= '1';
		radd1 <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '0');
		radd2 <= (0 => '1', 1 => '1', 2 => '0', 3 => '0', 4 => '0');
		wait for 100 ns;

    end process;

end architecture
